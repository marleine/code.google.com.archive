// FILE: Logic.vh

// ************************************************************************

// default verilog header file

// units of time and time resolution for this run
`timescale 1ps / 1ps

// this must be the very first module for interactive probing to work
module test;

// reg		a;
// wire		b;

// needed for interactive verilog probing.
   integer         tmp_channel;

// instantiate main verilog module
// NOTE: the name of the module must be the same as its type

	Logic Logic();

    initial
      begin
//    	$dumpfile();
//	$dumpvars;

//	a = 0;

// #1000 	a = 1; 

// #2000 	a = 0; 

//	$finish;
      end

endmodule

// include files
// `include "foo.v"

// ************************************************************************

// VERILOG netlist for "Logic" (generated by MMI_SUE4.4.0)

module xgate (in, in_L, t1, t2);
	inout		t1;
	inout		t2;
	input		in;
	input		in_L;
 
	pmos p(t2,t1,in_L);
	nmos n(t2,t1,in);

endmodule		// xgate

module my_xor (in1, in2, out);
	input		in1;
	input		in2;
	output		out;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	not #0 inv(net_1, in1);
	not #0 inv_1(out, net_2);
	not #0 inv_2(net_3, in2);
	xgate xgate(.in_L(net_1), .t2(net_2), .in(in1), .t1(in2));
	xgate xgate_1(.in(net_1), .t2(net_2), .t1(net_3), .in_L(in1));

endmodule		// my_xor

module MUX_2_1 (S0, a, b, out);
	input		S0;
	input		a;
	input		b;
	output		out;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	assign #0 net_1 = !(a && net_2);
	assign #0 net_3 = !(b && S0);
	assign #0 out = !(net_1 && net_3);
	not #0 inv(net_2, S0);

endmodule		// MUX_2_1

module MUX_4_1 (S, a, b, c, d, out);
	input		a;
	input		b;
	input		c;
	input		d;
	input	[1:0]	S;
	output		out;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	MUX_2_1 MUX_2_1(.S0(net_1), .out(net_2), .a(a), .b(b));
	MUX_2_1 MUX_2_2(.out(net_3), .b(d), .S0(S[0]), .a(c));
	MUX_2_1 MUX_2_3(.a(net_2), .b(net_3), .out(out), .S0(S[1]));
	not #0 inv(net_1, S[0]);

endmodule		// MUX_4_1

module Logic (Out, S, a, b);
	input		a;
	input		b;
	input	[1:0]	S;
	output		Out;
 
	wire		net_6;
	wire		net_2;
	wire		net_7;
	wire		net_3;
	wire		net_4;
	wire		net_5;
	wire		net_1;
 
	not #0 inv(net_5, net_6);
	not #0 inv_1(net_2, net_3);
	my_xor my_xor(.out(net_1), .in1(a), .in2(b));
	my_xor my_xor_1(.out(net_7), .in1(a), .in2(b));
	not #0 inv_2(net_4, net_7);
	assign #0 net_6 = !(a && b);
	assign net_3 = !(a || b);
	MUX_4_1 MUX_4_1(.c(net_1), .b(net_2), .d(net_4), .a(net_5), 
		.out(Out), .S(S[1:0]));

endmodule		// Logic

