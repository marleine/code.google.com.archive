// FILE: Comp.vh

// ************************************************************************

// default verilog header file

// units of time and time resolution for this run
`timescale 1ps / 1ps

// this must be the very first module for interactive probing to work
module test;

// reg		a;
// wire		b;

// needed for interactive verilog probing.
   integer         tmp_channel;

// instantiate main verilog module
// NOTE: the name of the module must be the same as its type

	Comp Comp();

    initial
      begin
//    	$dumpfile();
//	$dumpvars;

//	a = 0;

// #1000 	a = 1; 

// #2000 	a = 0; 

//	$finish;
      end

endmodule

// include files
// `include "foo.v"

// ************************************************************************

// VERILOG netlist for "Comp" (generated by MMI_SUE4.4.0)

module xgate (in, in_L, t1, t2);
	inout		t1;
	inout		t2;
	input		in;
	input		in_L;
 
	pmos p(t2,t1,in_L);
	nmos n(t2,t1,in);

endmodule		// xgate

module my_xor (in1, in2, out);
	input		in1;
	input		in2;
	output		out;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	not #0 inv(net_1, in1);
	not #0 inv_1(out, net_2);
	not #0 inv_2(net_3, in2);
	xgate xgate(.in_L(net_1), .t2(net_2), .in(in1), .t1(in2));
	xgate xgate_1(.in(net_1), .t2(net_2), .t1(net_3), .in_L(in1));

endmodule		// my_xor

module Comp (B, Out, S);
	input	[31:0]	B;
	input	[1:1]	S;
	output	[31:0]	Out;
 
	my_xor my_xor(.out(Out[31]), .in1(B[31]), .in2(S[1]));
	my_xor my_xor_1(.out(Out[30]), .in1(B[30]), .in2(S[1]));
	my_xor my_xor_2(.out(Out[29]), .in1(B[29]), .in2(S[1]));
	my_xor my_xor_3(.out(Out[28]), .in1(B[28]), .in2(S[1]));
	my_xor my_xor_4(.out(Out[27]), .in1(B[27]), .in2(S[1]));
	my_xor my_xor_5(.out(Out[26]), .in1(B[26]), .in2(S[1]));
	my_xor my_xor_6(.out(Out[25]), .in1(B[25]), .in2(S[1]));
	my_xor my_xor_7(.out(Out[24]), .in1(B[24]), .in2(S[1]));
	my_xor my_xor_8(.out(Out[23]), .in1(B[23]), .in2(S[1]));
	my_xor my_xor_9(.out(Out[22]), .in1(B[22]), .in2(S[1]));
	my_xor my_xor_10(.out(Out[21]), .in1(B[21]), .in2(S[1]));
	my_xor my_xor_11(.out(Out[20]), .in1(B[20]), .in2(S[1]));
	my_xor my_xor_12(.out(Out[19]), .in1(B[19]), .in2(S[1]));
	my_xor my_xor_13(.out(Out[18]), .in1(B[18]), .in2(S[1]));
	my_xor my_xor_14(.out(Out[17]), .in1(B[17]), .in2(S[1]));
	my_xor my_xor_15(.out(Out[16]), .in1(B[16]), .in2(S[1]));
	my_xor my_xor_16(.out(Out[15]), .in1(B[15]), .in2(S[1]));
	my_xor my_xor_17(.out(Out[14]), .in1(B[14]), .in2(S[1]));
	my_xor my_xor_18(.out(Out[13]), .in1(B[13]), .in2(S[1]));
	my_xor my_xor_19(.out(Out[12]), .in1(B[12]), .in2(S[1]));
	my_xor my_xor_20(.out(Out[11]), .in1(B[11]), .in2(S[1]));
	my_xor my_xor_21(.out(Out[10]), .in1(B[10]), .in2(S[1]));
	my_xor my_xor_22(.out(Out[9]), .in1(B[9]), .in2(S[1]));
	my_xor my_xor_23(.out(Out[8]), .in1(B[8]), .in2(S[1]));
	my_xor my_xor_24(.out(Out[7]), .in1(B[7]), .in2(S[1]));
	my_xor my_xor_25(.out(Out[6]), .in1(B[6]), .in2(S[1]));
	my_xor my_xor_26(.out(Out[5]), .in1(B[5]), .in2(S[1]));
	my_xor my_xor_27(.out(Out[4]), .in1(B[4]), .in2(S[1]));
	my_xor my_xor_28(.out(Out[3]), .in1(B[3]), .in2(S[1]));
	my_xor my_xor_29(.out(Out[2]), .in1(B[2]), .in2(S[1]));
	my_xor my_xor_30(.out(Out[1]), .in1(B[1]), .in2(S[1]));
	my_xor my_xor_31(.out(Out[0]), .in1(B[0]), .in2(S[1]));

endmodule		// Comp

