* FILE: Register_file_32bits.sp

********************** begin header *****************************

* Example header file for SPICE

.OPTIONS post ACCT OPTS lvltim=2
.OPTIONS post_version=9007

.option gmindc=   10.0p       

.options ADM_V_SUPPLY=3.3
*.options ADM_ACCURACY=10
*.options ADM_MODE=exp
.options ADM_MODE=acs
*.options ADM_MAXSTEP=10p
.options ignore_meas=0
*.param temper = 105

**################################################
* Corners are TT, SS, FF, SF, FS
.lib '<spice_model_file>' TT
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=2 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.35u
.param lp_min   =  0.35u

* used in source/drain area/perimeter calculation
.param sdd        =  0.95

.PARAM vddp=3.0		$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 10p 16n
*********************** end header ******************************

* SPICE netlist for "Register_file_32bits" (generated by MMI_SUE4.4.0)

.SUBCKT nand2 in0 in1 out WP=2 WN=2
M_1 out in0 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_2 out in0 net_1 gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_3 out in1 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_4 net_1 in1 gnd gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
.ENDS	$ nand2

.SUBCKT inverter in out WP=2 LP=lp_min WN=1 LN=ln_min
M_1 out in gnd gnd n W='WN*1u' L=LN ad='arean(WN,sdd)' as='arean(WN,sdd)' 
+ pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_2 out in vdd vdd p W='WP*1u' L=LP ad='areap(WP,sdd)' as='areap(WP,sdd)' 
+ pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
.ENDS	$ inverter

.SUBCKT writeEnable in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] 
+ in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] 
+ in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] 
+ in[29] in[30] in[31] out[0] out[1] out[2] out[3] out[4] out[5] out[6] 
+ out[7] out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15] 
+ out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23] out[24] 
+ out[25] out[26] out[27] out[28] out[29] out[30] out[31] writeBit 
Xnand2 in[0] writeBit net_31 nand2 
Xinverter net_31 out[0] inverter 
Xnand2_1 in[1] writeBit net_7 nand2 
Xinverter_1 net_7 out[1] inverter 
Xnand2_2 in[2] writeBit net_13 nand2 
Xinverter_2 net_13 out[2] inverter 
Xnand2_3 in[3] writeBit net_20 nand2 
Xinverter_3 net_20 out[3] inverter 
Xnand2_4 in[4] writeBit net_27 nand2 
Xinverter_4 net_27 out[4] inverter 
Xnand2_5 in[5] writeBit net_2 nand2 
Xinverter_5 net_2 out[5] inverter 
Xnand2_6 in[6] writeBit net_9 nand2 
Xinverter_6 net_9 out[6] inverter 
Xnand2_7 in[7] writeBit net_17 nand2 
Xinverter_7 net_17 out[7] inverter 
Xnand2_8 in[8] writeBit net_25 nand2 
Xinverter_8 net_25 out[8] inverter 
Xnand2_9 in[9] writeBit net_32 nand2 
Xinverter_9 net_32 out[9] inverter 
Xnand2_10 in[10] writeBit net_6 nand2 
Xinverter_10 net_6 out[10] inverter 
Xnand2_11 in[11] writeBit net_14 nand2 
Xinverter_11 net_14 out[11] inverter 
Xnand2_12 in[12] writeBit net_21 nand2 
Xinverter_12 net_21 out[12] inverter 
Xnand2_13 in[13] writeBit net_22 nand2 
Xinverter_13 net_22 out[13] inverter 
Xnand2_14 in[14] writeBit net_28 nand2 
Xinverter_14 net_28 out[14] inverter 
Xnand2_15 in[15] writeBit net_3 nand2 
Xinverter_15 net_3 out[15] inverter 
Xnand2_16 in[16] writeBit net_10 nand2 
Xinverter_16 net_10 out[16] inverter 
Xnand2_17 in[17] writeBit net_18 nand2 
Xinverter_17 net_18 out[17] inverter 
Xnand2_18 in[18] writeBit net_26 nand2 
Xinverter_18 net_26 out[18] inverter 
Xnand2_19 in[19] writeBit net_1 nand2 
Xinverter_19 net_1 out[19] inverter 
Xnand2_20 in[20] writeBit net_8 nand2 
Xinverter_20 net_8 out[20] inverter 
Xnand2_21 in[21] writeBit net_16 nand2 
Xinverter_21 net_16 out[21] inverter 
Xnand2_22 in[22] writeBit net_23 nand2 
Xinverter_22 net_23 out[22] inverter 
Xnand2_23 in[23] writeBit net_29 nand2 
Xinverter_23 net_29 out[23] inverter 
Xnand2_24 in[24] writeBit net_4 nand2 
Xinverter_24 net_4 out[24] inverter 
Xnand2_25 in[25] writeBit net_11 nand2 
Xinverter_25 net_11 out[25] inverter 
Xnand2_26 in[26] writeBit net_19 nand2 
Xinverter_26 net_19 out[26] inverter 
Xnand2_27 in[27] writeBit net_15 nand2 
Xinverter_27 net_15 out[27] inverter 
Xnand2_28 in[28] writeBit net_24 nand2 
Xinverter_28 net_24 out[28] inverter 
Xnand2_29 in[29] writeBit net_30 nand2 
Xinverter_29 net_30 out[29] inverter 
Xnand2_30 in[30] writeBit net_5 nand2 
Xinverter_30 net_5 out[30] inverter 
Xnand2_31 in[31] writeBit net_12 nand2 
Xinverter_31 net_12 out[31] inverter 
.ENDS	$ writeEnable

.SUBCKT nand3 in0 in1 in2 out WP=2 WN=3
M_1 out in0 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_2 out in0 net_1 gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_3 out in1 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_4 net_1 in1 net_2 gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_5 out in2 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_6 net_2 in2 gnd gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
.ENDS	$ nand3

.SUBCKT Dec_3x8 a[0] a[1] a[2] out2D[0] out2D[1] out2D[2] out2D[3] out2D[4] 
+ out2D[5] out2D[6] out2D[7] 
Xinverter a[0] net_1 inverter 
Xinverter_1 a[1] net_4 inverter 
Xinverter_2 a[2] net_2 inverter 
Xnand3 net_1 net_4 a[2] net_11 nand3 WN=2
Xinverter_3 net_11 out2D[1] inverter 
Xnand3_1 net_1 a[1] net_2 net_9 nand3 WN=2
Xinverter_4 net_9 out2D[2] inverter 
Xnand3_2 net_1 a[1] a[2] net_6 nand3 WN=2
Xinverter_5 net_6 out2D[3] inverter 
Xnand3_3 a[0] net_4 net_2 net_10 nand3 WN=2
Xinverter_6 net_10 out2D[4] inverter 
Xnand3_4 a[0] net_4 a[2] net_8 nand3 WN=2
Xinverter_7 net_8 out2D[5] inverter 
Xnand3_5 a[0] a[1] net_2 net_3 nand3 WN=2
Xinverter_8 net_3 out2D[6] inverter 
Xnand3_6 a[0] a[1] a[2] net_5 nand3 WN=2
Xinverter_9 net_5 out2D[7] inverter 
Xnand3_7 net_1 net_4 net_2 net_7 nand3 WN=2
Xinverter_10 net_7 out2D[0] inverter 
.ENDS	$ Dec_3x8

.SUBCKT Dec_2x4 a[0] a[1] enable outD[0] outD[1] outD[2] outD[3] 
Xinverter a[0] net_4 inverter 
Xinverter_1 a[1] net_2 inverter 
Xnand3 enable net_4 net_2 net_8 nand3 WN=2
Xinverter_2 a[1] net_1 inverter 
Xnand3_1 enable a[0] net_1 net_7 nand3 WN=2
Xnand3_2 enable net_5 a[1] net_6 nand3 WN=2
Xinverter_3 a[0] net_5 inverter 
Xnand3_3 enable a[0] a[1] net_3 nand3 WN=2
Xinverter_4 net_8 outD[0] inverter 
Xinverter_5 net_7 outD[1] inverter 
Xinverter_6 net_6 outD[2] inverter 
Xinverter_7 net_3 outD[3] inverter 
.ENDS	$ Dec_2x4

.SUBCKT Dec_5x32 in[0] in[1] in[2] in[3] in[4] outD5[0] outD5[1] outD5[2] 
+ outD5[3] outD5[4] outD5[5] outD5[6] outD5[7] outD5[8] outD5[9] outD5[10] 
+ outD5[11] outD5[12] outD5[13] outD5[14] outD5[15] outD5[16] outD5[17] 
+ outD5[18] outD5[19] outD5[20] outD5[21] outD5[22] outD5[23] outD5[24] 
+ outD5[25] outD5[26] outD5[27] outD5[28] outD5[29] outD5[30] outD5[31] 
XDec_3x8 in[2] in[3] in[4] out[0] out[1] out[2] out[3] out[4] out[5] out[6] 
+ out[7] Dec_3x8 
XDec_2x4 in[0] in[1] out[0] outD5[0] outD5[1] outD5[2] outD5[3] Dec_2x4 
XDec_2x4_1 in[0] in[1] out[1] outD5[4] outD5[5] outD5[6] outD5[7] Dec_2x4 
XDec_2x4_2 in[0] in[1] out[2] outD5[8] outD5[9] outD5[10] outD5[11] Dec_2x4 
+ 
XDec_2x4_3 in[0] in[1] out[3] outD5[12] outD5[13] outD5[14] outD5[15] 
+ Dec_2x4 
XDec_2x4_4 in[0] in[1] out[4] outD5[16] outD5[17] outD5[18] outD5[19] 
+ Dec_2x4 
XDec_2x4_5 in[0] in[1] out[5] outD5[20] outD5[21] outD5[22] outD5[23] 
+ Dec_2x4 
XDec_2x4_6 in[0] in[1] out[6] outD5[24] outD5[25] outD5[26] outD5[27] 
+ Dec_2x4 
XDec_2x4_7 in[0] in[1] out[7] outD5[28] outD5[29] outD5[30] outD5[31] 
+ Dec_2x4 
.ENDS	$ Dec_5x32

.SUBCKT Reg0_1bit R1 R2 out1 out2 
M_1 out1 R1 gnd gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' as='arean(1,sdd)' 
+ pd='perin(1,sdd)' ps='perin(1,sdd)' 
M_2 out2 R2 gnd gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' as='arean(1,sdd)' 
+ pd='perin(1,sdd)' ps='perin(1,sdd)' 
.ENDS	$ Reg0_1bit

.SUBCKT Reg0_32bit R1 R2 out1[0] out1[1] out1[2] out1[3] out1[4] out1[5] 
+ out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] out1[13] 
+ out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] out1[21] 
+ out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] out1[29] 
+ out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] out2[5] out2[6] 
+ out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] out2[13] out2[14] 
+ out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] out2[21] out2[22] 
+ out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] out2[29] out2[30] 
+ out2[31] 
XReg0_1bit R1 R2 out1[0] out2[0] Reg0_1bit 
XReg0_1bit_1 R1 R2 out1[1] out2[1] Reg0_1bit 
XReg0_1bit_2 R1 R2 out1[2] out2[2] Reg0_1bit 
XReg0_1bit_3 R1 R2 out1[3] out2[3] Reg0_1bit 
XReg0_1bit_4 R1 R2 out1[4] out2[4] Reg0_1bit 
XReg0_1bit_5 R1 R2 out1[5] out2[5] Reg0_1bit 
XReg0_1bit_6 R1 R2 out1[6] out2[6] Reg0_1bit 
XReg0_1bit_7 R1 R2 out1[7] out2[7] Reg0_1bit 
XReg0_1bit_8 R1 R2 out1[8] out2[8] Reg0_1bit 
XReg0_1bit_9 R1 R2 out1[9] out2[9] Reg0_1bit 
XReg0_1bit_10 R1 R2 out1[10] out2[10] Reg0_1bit 
XReg0_1bit_11 R1 R2 out1[11] out2[11] Reg0_1bit 
XReg0_1bit_12 R1 R2 out1[12] out2[12] Reg0_1bit 
XReg0_1bit_13 R1 R2 out1[13] out2[13] Reg0_1bit 
XReg0_1bit_14 R1 R2 out1[14] out2[14] Reg0_1bit 
XReg0_1bit_15 R1 R2 out1[15] out2[15] Reg0_1bit 
XReg0_1bit_16 R1 R2 out1[16] out2[16] Reg0_1bit 
XReg0_1bit_17 R1 R2 out1[17] out2[17] Reg0_1bit 
XReg0_1bit_18 R1 R2 out1[18] out2[18] Reg0_1bit 
XReg0_1bit_19 R1 R2 out1[19] out2[19] Reg0_1bit 
XReg0_1bit_20 R1 R2 out1[20] out2[20] Reg0_1bit 
XReg0_1bit_21 R1 R2 out1[21] out2[21] Reg0_1bit 
XReg0_1bit_22 R1 R2 out1[22] out2[22] Reg0_1bit 
XReg0_1bit_23 R1 R2 out1[23] out2[23] Reg0_1bit 
XReg0_1bit_24 R1 R2 out1[24] out2[24] Reg0_1bit 
XReg0_1bit_25 R1 R2 out1[25] out2[25] Reg0_1bit 
XReg0_1bit_26 R1 R2 out1[26] out2[26] Reg0_1bit 
XReg0_1bit_27 R1 R2 out1[27] out2[27] Reg0_1bit 
XReg0_1bit_28 R1 R2 out1[28] out2[28] Reg0_1bit 
XReg0_1bit_29 R1 R2 out1[29] out2[29] Reg0_1bit 
XReg0_1bit_30 R1 R2 out1[30] out2[30] Reg0_1bit 
XReg0_1bit_31 R1 R2 out1[31] out2[31] Reg0_1bit 
.ENDS	$ Reg0_32bit

.SUBCKT Reg_1bit R1 R2 data out1 out2 write 
Xinverter net_2 net_1 inverter 
M_1 net_1 write net_3 gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' 
+ as='arean(1,sdd)' pd='perin(1,sdd)' ps='perin(1,sdd)' M=4
Xinverter_1 net_1 net_2 inverter M=4
Xinverter_2 data net_3 inverter M=4
M_2 out1 R1 net_2 gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' 
+ as='arean(1,sdd)' pd='perin(1,sdd)' ps='perin(1,sdd)' 
M_3 out2 R2 net_2 gnd n W='1*1u' L=ln_min ad='arean(1,sdd)' 
+ as='arean(1,sdd)' pd='perin(1,sdd)' ps='perin(1,sdd)' 
.ENDS	$ Reg_1bit

.SUBCKT Reg_32bit R1 R2 data[0] data[1] data[2] data[3] data[4] data[5] 
+ data[6] data[7] data[8] data[9] data[10] data[11] data[12] data[13] 
+ data[14] data[15] data[16] data[17] data[18] data[19] data[20] data[21] 
+ data[22] data[23] data[24] data[25] data[26] data[27] data[28] data[29] 
+ data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] out1[5] out1[6] 
+ out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] out1[13] out1[14] 
+ out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] out1[21] out1[22] 
+ out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] out1[29] out1[30] 
+ out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] out2[5] out2[6] out2[7] 
+ out2[8] out2[9] out2[10] out2[11] out2[12] out2[13] out2[14] out2[15] 
+ out2[16] out2[17] out2[18] out2[19] out2[20] out2[21] out2[22] out2[23] 
+ out2[24] out2[25] out2[26] out2[27] out2[28] out2[29] out2[30] out2[31] 
+ write 
XReg_1bit R1 R2 data[0] out1[0] out2[0] write Reg_1bit 
XReg_1bit_1 R1 R2 data[1] out1[1] out2[1] write Reg_1bit 
XReg_1bit_2 R1 R2 data[2] out1[2] out2[2] write Reg_1bit 
XReg_1bit_3 R1 R2 data[3] out1[3] out2[3] write Reg_1bit 
XReg_1bit_4 R1 R2 data[4] out1[4] out2[4] write Reg_1bit 
XReg_1bit_5 R1 R2 data[5] out1[5] out2[5] write Reg_1bit 
XReg_1bit_6 R1 R2 data[6] out1[6] out2[6] write Reg_1bit 
XReg_1bit_7 R1 R2 data[7] out1[7] out2[7] write Reg_1bit 
XReg_1bit_8 R1 R2 data[8] out1[8] out2[8] write Reg_1bit 
XReg_1bit_9 R1 R2 data[9] out1[9] out2[9] write Reg_1bit 
XReg_1bit_10 R1 R2 data[10] out1[10] out2[10] write Reg_1bit 
XReg_1bit_11 R1 R2 data[11] out1[11] out2[11] write Reg_1bit 
XReg_1bit_12 R1 R2 data[12] out1[12] out2[12] write Reg_1bit 
XReg_1bit_13 R1 R2 data[13] out1[13] out2[13] write Reg_1bit 
XReg_1bit_14 R1 R2 data[14] out1[14] out2[14] write Reg_1bit 
XReg_1bit_15 R1 R2 data[15] out1[15] out2[15] write Reg_1bit 
XReg_1bit_16 R1 R2 data[16] out1[16] out2[16] write Reg_1bit 
XReg_1bit_17 R1 R2 data[17] out1[17] out2[17] write Reg_1bit 
XReg_1bit_18 R1 R2 data[18] out1[18] out2[18] write Reg_1bit 
XReg_1bit_19 R1 R2 data[19] out1[19] out2[19] write Reg_1bit 
XReg_1bit_20 R1 R2 data[20] out1[20] out2[20] write Reg_1bit 
XReg_1bit_21 R1 R2 data[21] out1[21] out2[21] write Reg_1bit 
XReg_1bit_22 R1 R2 data[22] out1[22] out2[22] write Reg_1bit 
XReg_1bit_23 R1 R2 data[23] out1[23] out2[23] write Reg_1bit 
XReg_1bit_24 R1 R2 data[24] out1[24] out2[24] write Reg_1bit 
XReg_1bit_25 R1 R2 data[25] out1[25] out2[25] write Reg_1bit 
XReg_1bit_26 R1 R2 data[26] out1[26] out2[26] write Reg_1bit 
XReg_1bit_27 R1 R2 data[27] out1[27] out2[27] write Reg_1bit 
XReg_1bit_28 R1 R2 data[28] out1[28] out2[28] write Reg_1bit 
XReg_1bit_29 R1 R2 data[29] out1[29] out2[29] write Reg_1bit 
XReg_1bit_30 R1 R2 data[30] out1[30] out2[30] write Reg_1bit 
XReg_1bit_31 R1 R2 data[31] out1[31] out2[31] write Reg_1bit 
.ENDS	$ Reg_32bit

* start main CELL Register_file_32bits
* .SUBCKT Register_file_32bits address_read1[0] address_read1[1] 
*+ address_read1[2] address_read1[3] address_read1[4] address_read2[0] 
*+ address_read2[1] address_read2[2] address_read2[3] address_read2[4] 
*+ address_write[0] address_write[1] address_write[2] address_write[3] 
*+ address_write[4] data[0] data[1] data[2] data[3] data[4] data[5] data[6] 
*+ data[7] data[8] data[9] data[10] data[11] data[12] data[13] data[14] 
*+ data[15] data[16] data[17] data[18] data[19] data[20] data[21] data[22] 
*+ data[23] data[24] data[25] data[26] data[27] data[28] data[29] data[30] 
*+ data[31] out1[0] out1[1] out1[2] out1[3] out1[4] out1[5] out1[6] out1[7] 
*+ out1[8] out1[9] out1[10] out1[11] out1[12] out1[13] out1[14] out1[15] 
*+ out1[16] out1[17] out1[18] out1[19] out1[20] out1[21] out1[22] out1[23] 
*+ out1[24] out1[25] out1[26] out1[27] out1[28] out1[29] out1[30] out1[31] 
*+ out2[0] out2[1] out2[2] out2[3] out2[4] out2[5] out2[6] out2[7] out2[8] 
*+ out2[9] out2[10] out2[11] out2[12] out2[13] out2[14] out2[15] out2[16] 
*+ out2[17] out2[18] out2[19] out2[20] out2[21] out2[22] out2[23] out2[24] 
*+ out2[25] out2[26] out2[27] out2[28] out2[29] out2[30] out2[31] 
*+ write_enable 
XwriteEnable net_1[0] net_1[1] net_1[2] net_1[3] net_1[4] net_1[5] net_1[6] 
+ net_1[7] net_1[8] net_1[9] net_1[10] net_1[11] net_1[12] net_1[13] 
+ net_1[14] net_1[15] net_1[16] net_1[17] net_1[18] net_1[19] net_1[20] 
+ net_1[21] net_1[22] net_1[23] net_1[24] net_1[25] net_1[26] net_1[27] 
+ net_1[28] net_1[29] net_1[30] net_1[31] w[0] w[1] w[2] w[3] w[4] w[5] 
+ w[6] w[7] w[8] w[9] w[10] w[11] w[12] w[13] w[14] w[15] w[16] w[17] w[18] 
+ w[19] w[20] w[21] w[22] w[23] w[24] w[25] w[26] w[27] w[28] w[29] w[30] 
+ w[31] write_enable writeEnable 
XDec_5x32 address_write[0] address_write[1] address_write[2] 
+ address_write[3] address_write[4] net_1[0] net_1[1] net_1[2] net_1[3] 
+ net_1[4] net_1[5] net_1[6] net_1[7] net_1[8] net_1[9] net_1[10] net_1[11] 
+ net_1[12] net_1[13] net_1[14] net_1[15] net_1[16] net_1[17] net_1[18] 
+ net_1[19] net_1[20] net_1[21] net_1[22] net_1[23] net_1[24] net_1[25] 
+ net_1[26] net_1[27] net_1[28] net_1[29] net_1[30] net_1[31] Dec_5x32 
XDec_5x32_1 address_read2[0] address_read2[1] address_read2[2] 
+ address_read2[3] address_read2[4] R2[0] R2[1] R2[2] R2[3] R2[4] R2[5] 
+ R2[6] R2[7] R2[8] R2[9] R2[10] R2[11] R2[12] R2[13] R2[14] R2[15] R2[16] 
+ R2[17] R2[18] R2[19] R2[20] R2[21] R2[22] R2[23] R2[24] R2[25] R2[26] 
+ R2[27] R2[28] R2[29] R2[30] R2[31] Dec_5x32 
XDec_5x32_2 address_read1[0] address_read1[1] address_read1[2] 
+ address_read1[3] address_read1[4] R1[0] R1[1] R1[2] R1[3] R1[4] R1[5] 
+ R1[6] R1[7] R1[8] R1[9] R1[10] R1[11] R1[12] R1[13] R1[14] R1[15] R1[16] 
+ R1[17] R1[18] R1[19] R1[20] R1[21] R1[22] R1[23] R1[24] R1[25] R1[26] 
+ R1[27] R1[28] R1[29] R1[30] R1[31] Dec_5x32 
XReg0_32bit inR1[0] inR2[0] out1[0] out1[1] out1[2] out1[3] out1[4] out1[5] 
+ out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] out1[13] 
+ out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] out1[21] 
+ out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] out1[29] 
+ out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] out2[5] out2[6] 
+ out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] out2[13] out2[14] 
+ out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] out2[21] out2[22] 
+ out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] out2[29] out2[30] 
+ out2[31] Reg0_32bit 
XReg_32bit inR1[1] inR2[1] data[0] data[1] data[2] data[3] data[4] data[5] 
+ data[6] data[7] data[8] data[9] data[10] data[11] data[12] data[13] 
+ data[14] data[15] data[16] data[17] data[18] data[19] data[20] data[21] 
+ data[22] data[23] data[24] data[25] data[26] data[27] data[28] data[29] 
+ data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] out1[5] out1[6] 
+ out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] out1[13] out1[14] 
+ out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] out1[21] out1[22] 
+ out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] out1[29] out1[30] 
+ out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] out2[5] out2[6] out2[7] 
+ out2[8] out2[9] out2[10] out2[11] out2[12] out2[13] out2[14] out2[15] 
+ out2[16] out2[17] out2[18] out2[19] out2[20] out2[21] out2[22] out2[23] 
+ out2[24] out2[25] out2[26] out2[27] out2[28] out2[29] out2[30] out2[31] 
+ w[1] Reg_32bit 
XReg_32bit_1 inR1[2] inR2[2] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[2] Reg_32bit 
XReg_32bit_2 inR1[3] inR2[3] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[3] Reg_32bit 
XReg_32bit_3 inR1[4] inR2[4] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[4] Reg_32bit 
XReg_32bit_4 inR1[5] inR2[5] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[5] Reg_32bit 
XReg_32bit_5 inR1[6] inR2[6] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[6] Reg_32bit 
XReg_32bit_6 inR1[7] inR2[7] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[7] Reg_32bit 
XReg_32bit_7 inR1[8] inR2[8] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[8] Reg_32bit 
XReg_32bit_8 inR1[9] inR2[9] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[9] Reg_32bit 
XReg_32bit_9 inR1[10] inR2[10] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[10] Reg_32bit 
XReg_32bit_10 inR1[11] inR2[11] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[11] Reg_32bit 
XReg_32bit_11 inR1[12] inR2[12] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[12] Reg_32bit 
XReg_32bit_12 inR1[13] inR2[13] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[13] Reg_32bit 
XReg_32bit_13 inR1[14] inR2[14] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[14] Reg_32bit 
XReg_32bit_14 inR1[15] inR2[15] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[15] Reg_32bit 
XReg_32bit_15 inR1[16] inR2[16] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[16] Reg_32bit 
XReg_32bit_16 inR1[17] inR2[17] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[17] Reg_32bit 
XReg_32bit_17 inR1[18] inR2[18] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[18] Reg_32bit 
XReg_32bit_18 inR1[19] inR2[19] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[19] Reg_32bit 
XReg_32bit_19 inR1[20] inR2[20] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[20] Reg_32bit 
XReg_32bit_20 inR1[21] inR2[21] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[21] Reg_32bit 
XReg_32bit_21 inR1[22] inR2[22] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[22] Reg_32bit 
XReg_32bit_22 inR1[23] inR2[23] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[23] Reg_32bit 
XReg_32bit_23 inR1[24] inR2[24] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[24] Reg_32bit 
XReg_32bit_24 inR1[25] inR2[25] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[25] Reg_32bit 
XReg_32bit_25 inR1[26] inR2[26] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[26] Reg_32bit 
XReg_32bit_26 inR1[27] inR2[27] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[27] Reg_32bit 
XReg_32bit_27 inR1[28] inR2[28] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[28] Reg_32bit 
XReg_32bit_28 inR1[29] inR2[29] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[29] Reg_32bit 
XReg_32bit_29 inR1[30] inR2[30] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[30] Reg_32bit 
XReg_32bit_30 inR1[31] inR2[31] data[0] data[1] data[2] data[3] data[4] 
+ data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] 
+ data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] 
+ data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] 
+ data[29] data[30] data[31] out1[0] out1[1] out1[2] out1[3] out1[4] 
+ out1[5] out1[6] out1[7] out1[8] out1[9] out1[10] out1[11] out1[12] 
+ out1[13] out1[14] out1[15] out1[16] out1[17] out1[18] out1[19] out1[20] 
+ out1[21] out1[22] out1[23] out1[24] out1[25] out1[26] out1[27] out1[28] 
+ out1[29] out1[30] out1[31] out2[0] out2[1] out2[2] out2[3] out2[4] 
+ out2[5] out2[6] out2[7] out2[8] out2[9] out2[10] out2[11] out2[12] 
+ out2[13] out2[14] out2[15] out2[16] out2[17] out2[18] out2[19] out2[20] 
+ out2[21] out2[22] out2[23] out2[24] out2[25] out2[26] out2[27] out2[28] 
+ out2[29] out2[30] out2[31] w[31] Reg_32bit 
* .ENDS	$ Register_file_32bits

.GLOBAL gnd vdd

.END

