* FILE: MUX_64_32.sp

********************** begin header *****************************

* Example header file for SPICE

.OPTIONS post ACCT OPTS lvltim=2
.OPTIONS post_version=9007

.option gmindc=   10.0p       

.options ADM_V_SUPPLY=3.3
*.options ADM_ACCURACY=10
*.options ADM_MODE=exp
.options ADM_MODE=acs
*.options ADM_MAXSTEP=10p
.options ignore_meas=0
*.param temper = 105

**################################################
* Corners are TT, SS, FF, SF, FS
.lib '<spice_model_file>' TT
**################################################

.param  arean(w,sdd) = '(w*sdd*1p)'
.param  areap(w,sdd) = '(w*sdd*1p)'
* Setup either one or the other of the following
* For ACM=2 fet models
.param  perin(w,sdd) = '(2u*(w+sdd))'
.param  perip(w,sdd) = '(2u*(w+sdd))'
* For ACM=3 fet models
*.param  perin(w,sdd) = '(1u*(w+2*sdd))'
*.param  perip(w,sdd) = '(1u*(w+2*sdd))'

.param ln_min   =  0.35u
.param lp_min   =  0.35u

* used in source/drain area/perimeter calculation
.param sdd        =  0.95

.PARAM vddp=3.0		$ VDD voltage

VDD vdd 0 DC vddp 

.TEMP 105
.TRAN 10p 16n
*********************** end header ******************************

* SPICE netlist for "MUX_64_32" (generated by MMI_SUE4.4.0)

.SUBCKT nand2 in0 in1 out WP=2 WN=2
M_1 out in0 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_2 out in0 net_1 gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_3 out in1 vdd vdd p W='WP*1u' L=lp_min ad='areap(WP,sdd)' 
+ as='areap(WP,sdd)' pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
M_4 net_1 in1 gnd gnd n W='WN*1u' L=ln_min ad='arean(WN,sdd)' 
+ as='arean(WN,sdd)' pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
.ENDS	$ nand2

.SUBCKT inverter in out WP=2 LP=lp_min WN=1 LN=ln_min
M_1 out in gnd gnd n W='WN*1u' L=LN ad='arean(WN,sdd)' as='arean(WN,sdd)' 
+ pd='perin(WN,sdd)' ps='perin(WN,sdd)' 
M_2 out in vdd vdd p W='WP*1u' L=LP ad='areap(WP,sdd)' as='areap(WP,sdd)' 
+ pd='perip(WP,sdd)' ps='perip(WP,sdd)' 
.ENDS	$ inverter

.SUBCKT MUX_2_1 S0 a b out 
Xnand2 a net_1 net_2 nand2 
Xnand2_1 b S0 net_3 nand2 
Xnand2_2 net_2 net_3 out nand2 
Xinverter S0 net_1 inverter 
.ENDS	$ MUX_2_1

* start main CELL MUX_64_32
* .SUBCKT MUX_64_32 A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] A[8] A[9] A[10] 
*+ A[11] A[12] A[13] A[14] A[15] A[16] A[17] A[18] A[19] A[20] A[21] A[22] 
*+ A[23] A[24] A[25] A[26] A[27] A[28] A[29] A[30] A[31] B[0] B[1] B[2] 
*+ B[3] B[4] B[5] B[6] B[7] B[8] B[9] B[10] B[11] B[12] B[13] B[14] B[15] 
*+ B[16] B[17] B[18] B[19] B[20] B[21] B[22] B[23] B[24] B[25] B[26] B[27] 
*+ B[28] B[29] B[30] B[31] Out[0] Out[1] Out[2] Out[3] Out[4] Out[5] Out[6] 
*+ Out[7] Out[8] Out[9] Out[10] Out[11] Out[12] Out[13] Out[14] Out[15] 
*+ Out[16] Out[17] Out[18] Out[19] Out[20] Out[21] Out[22] Out[23] Out[24] 
*+ Out[25] Out[26] Out[27] Out[28] Out[29] Out[30] Out[31] S[2] 
XMUX_2_1 S[2] A[0] B[0] Out[0] MUX_2_1 
XMUX_2_2 S[2] A[1] B[1] Out[1] MUX_2_1 
XMUX_2_3 S[2] A[2] B[2] Out[2] MUX_2_1 
XMUX_2_4 S[2] A[3] B[3] Out[3] MUX_2_1 
XMUX_2_5 S[2] A[4] B[4] Out[4] MUX_2_1 
XMUX_2_6 S[2] A[5] B[5] Out[5] MUX_2_1 
XMUX_2_7 S[2] A[6] B[6] Out[6] MUX_2_1 
XMUX_2_8 S[2] A[7] B[7] Out[7] MUX_2_1 
XMUX_2_9 S[2] A[8] B[8] Out[8] MUX_2_1 
XMUX_2_10 S[2] A[9] B[9] Out[9] MUX_2_1 
XMUX_2_11 S[2] A[10] B[10] Out[10] MUX_2_1 
XMUX_2_12 S[2] A[11] B[11] Out[11] MUX_2_1 
XMUX_2_13 S[2] A[12] B[12] Out[12] MUX_2_1 
XMUX_2_14 S[2] A[13] B[13] Out[13] MUX_2_1 
XMUX_2_15 S[2] A[14] B[14] Out[14] MUX_2_1 
XMUX_2_16 S[2] A[15] B[15] Out[15] MUX_2_1 
XMUX_2_17 S[2] A[16] B[16] Out[16] MUX_2_1 
XMUX_2_18 S[2] A[17] B[17] Out[17] MUX_2_1 
XMUX_2_19 S[2] A[18] B[18] Out[18] MUX_2_1 
XMUX_2_20 S[2] A[19] B[19] Out[19] MUX_2_1 
XMUX_2_21 S[2] A[20] B[20] Out[20] MUX_2_1 
XMUX_2_22 S[2] A[21] B[21] Out[21] MUX_2_1 
XMUX_2_23 S[2] A[22] B[22] Out[22] MUX_2_1 
XMUX_2_24 S[2] A[23] B[23] Out[23] MUX_2_1 
XMUX_2_25 S[2] A[24] B[24] Out[24] MUX_2_1 
XMUX_2_26 S[2] A[25] B[25] Out[25] MUX_2_1 
XMUX_2_27 S[2] A[26] B[26] Out[26] MUX_2_1 
XMUX_2_28 S[2] A[27] B[27] Out[27] MUX_2_1 
XMUX_2_29 S[2] A[28] B[28] Out[28] MUX_2_1 
XMUX_2_30 S[2] A[29] B[29] Out[29] MUX_2_1 
XMUX_2_31 S[2] A[30] B[30] Out[30] MUX_2_1 
XMUX_2_32 S[2] A[31] B[31] Out[31] MUX_2_1 
* .ENDS	$ MUX_64_32

.GLOBAL gnd vdd

.END

