// FILE: MUX_64_32.vh

// ************************************************************************

// default verilog header file

// units of time and time resolution for this run
`timescale 1ps / 1ps

// this must be the very first module for interactive probing to work
module test;

// reg		a;
// wire		b;

// needed for interactive verilog probing.
   integer         tmp_channel;

// instantiate main verilog module
// NOTE: the name of the module must be the same as its type

	MUX_64_32 MUX_64_32();

    initial
      begin
//    	$dumpfile();
//	$dumpvars;

//	a = 0;

// #1000 	a = 1; 

// #2000 	a = 0; 

//	$finish;
      end

endmodule

// include files
// `include "foo.v"

// ************************************************************************

// VERILOG netlist for "MUX_64_32" (generated by MMI_SUE4.4.0)

module MUX_2_1 (S0, a, b, out);
	input		S0;
	input		a;
	input		b;
	output		out;
 
	wire		net_2;
	wire		net_3;
	wire		net_1;
 
	assign #0 net_1 = !(a && net_2);
	assign #0 net_3 = !(b && S0);
	assign #0 out = !(net_1 && net_3);
	not #0 inv(net_2, S0);

endmodule		// MUX_2_1

module MUX_64_32 (A, B, Out, S);
	input	[31:0]	A;
	input	[31:0]	B;
	input	[2:2]	S;
	output	[31:0]	Out;
 
	MUX_2_1 MUX_2_1(.out(Out[0]), .a(A[0]), .b(B[0]), .S0(S[2]));
	MUX_2_1 MUX_2_2(.out(Out[1]), .a(A[1]), .b(B[1]), .S0(S[2]));
	MUX_2_1 MUX_2_3(.out(Out[2]), .a(A[2]), .b(B[2]), .S0(S[2]));
	MUX_2_1 MUX_2_4(.out(Out[3]), .a(A[3]), .b(B[3]), .S0(S[2]));
	MUX_2_1 MUX_2_5(.out(Out[4]), .a(A[4]), .b(B[4]), .S0(S[2]));
	MUX_2_1 MUX_2_6(.out(Out[5]), .a(A[5]), .b(B[5]), .S0(S[2]));
	MUX_2_1 MUX_2_7(.out(Out[6]), .a(A[6]), .b(B[6]), .S0(S[2]));
	MUX_2_1 MUX_2_8(.out(Out[7]), .a(A[7]), .b(B[7]), .S0(S[2]));
	MUX_2_1 MUX_2_9(.out(Out[8]), .a(A[8]), .b(B[8]), .S0(S[2]));
	MUX_2_1 MUX_2_10(.out(Out[9]), .a(A[9]), .b(B[9]), .S0(S[2]));
	MUX_2_1 MUX_2_11(.out(Out[10]), .a(A[10]), .b(B[10]), .S0(S[2]));
	MUX_2_1 MUX_2_12(.out(Out[11]), .a(A[11]), .b(B[11]), .S0(S[2]));
	MUX_2_1 MUX_2_13(.out(Out[12]), .a(A[12]), .b(B[12]), .S0(S[2]));
	MUX_2_1 MUX_2_14(.out(Out[13]), .a(A[13]), .b(B[13]), .S0(S[2]));
	MUX_2_1 MUX_2_15(.out(Out[14]), .a(A[14]), .b(B[14]), .S0(S[2]));
	MUX_2_1 MUX_2_16(.out(Out[15]), .a(A[15]), .b(B[15]), .S0(S[2]));
	MUX_2_1 MUX_2_17(.out(Out[16]), .a(A[16]), .b(B[16]), .S0(S[2]));
	MUX_2_1 MUX_2_18(.out(Out[17]), .a(A[17]), .b(B[17]), .S0(S[2]));
	MUX_2_1 MUX_2_19(.out(Out[18]), .a(A[18]), .b(B[18]), .S0(S[2]));
	MUX_2_1 MUX_2_20(.out(Out[19]), .a(A[19]), .b(B[19]), .S0(S[2]));
	MUX_2_1 MUX_2_21(.out(Out[20]), .a(A[20]), .b(B[20]), .S0(S[2]));
	MUX_2_1 MUX_2_22(.out(Out[21]), .a(A[21]), .b(B[21]), .S0(S[2]));
	MUX_2_1 MUX_2_23(.out(Out[22]), .a(A[22]), .b(B[22]), .S0(S[2]));
	MUX_2_1 MUX_2_24(.out(Out[23]), .a(A[23]), .b(B[23]), .S0(S[2]));
	MUX_2_1 MUX_2_25(.out(Out[24]), .a(A[24]), .b(B[24]), .S0(S[2]));
	MUX_2_1 MUX_2_26(.out(Out[25]), .a(A[25]), .b(B[25]), .S0(S[2]));
	MUX_2_1 MUX_2_27(.out(Out[26]), .a(A[26]), .b(B[26]), .S0(S[2]));
	MUX_2_1 MUX_2_28(.out(Out[27]), .a(A[27]), .b(B[27]), .S0(S[2]));
	MUX_2_1 MUX_2_29(.out(Out[28]), .a(A[28]), .b(B[28]), .S0(S[2]));
	MUX_2_1 MUX_2_30(.out(Out[29]), .a(A[29]), .b(B[29]), .S0(S[2]));
	MUX_2_1 MUX_2_31(.out(Out[30]), .a(A[30]), .b(B[30]), .S0(S[2]));
	MUX_2_1 MUX_2_32(.out(Out[31]), .a(A[31]), .b(B[31]), .S0(S[2]));

endmodule		// MUX_64_32

